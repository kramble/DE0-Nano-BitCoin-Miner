// Testbench for fpgaminer_top.v
// Assumes 50MHz clock and 500kbps comms, so bit period is 100 clock cycles

`timescale 1ns/1ps

module test_serial_icarus2();

	reg clk = 1'b0;
	reg RxD = 1'b1;	// Active low
	wire TxD;
	// wire led_out;
	wire led1, led2, led3;
	
	fpgaminer_top #(.SIM_SERIAL(1),.NUM_HASHERS(6),.LOOP(11),.SPEED_MHZ(50),.ICARUS(1)) uut 
		(clk, RxD, TxD, led1, led2, led3);
	
	reg [31:0] cycle = 32'd0;

	initial begin
		clk = 0;

		#100

		// Not setting uut.nonce as icarus protocol resets nonce on loading work
		// Aiming for match at t~44,000,000nS (it takes that long to count up from zero) - hashers 3
		// Aiming for match at t~25,000,000nS (it takes that long to count up from zero) - hashers 6
		
		while(1)
		begin
			#5 clk = 1; #5 clk = 0;

			// cgminer icarus detect ...
			// uut.midstate_buf = 256'h4679ba4ec99876bf4bfe086082b400254df6c356451471139a3afa71e48f544a;
			// uut.data_buf = 512'h0000028000000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000087320b1a1426674f2fa722ce;
			// uut.nonce = 32'h00018790;	// For 32'h000187a2

			// This is ever so crude (should be possible in verilog, but I wrote C code to generate it)
            // Send 4679ba4ec99876bf4bfe086082b400254df6c356451471139a3afa71e48f544a 0000000000000000000000000000000000000000 87320b1a1426674f2fa722ce

			// 100 clock cycle bit period, 8 bit, no parity, one start, 8 bits LSB first, one stop, 1=high

if(cycle==200)RxD<=0;
if(cycle==300)RxD<=0;
if(cycle==400)RxD<=1;
if(cycle==500)RxD<=1;
if(cycle==600)RxD<=0;
if(cycle==700)RxD<=0;
if(cycle==800)RxD<=0;
if(cycle==900)RxD<=1;
if(cycle==1000)RxD<=0;
if(cycle==1100)RxD<=1;
if(cycle==1200)RxD<=0;
if(cycle==1300)RxD<=1;
if(cycle==1400)RxD<=0;
if(cycle==1500)RxD<=0;
if(cycle==1600)RxD<=1;
if(cycle==1700)RxD<=1;
if(cycle==1800)RxD<=1;
if(cycle==1900)RxD<=1;
if(cycle==2000)RxD<=0;
if(cycle==2100)RxD<=1;
if(cycle==2200)RxD<=0;
if(cycle==2300)RxD<=0;
if(cycle==2400)RxD<=1;
if(cycle==2500)RxD<=0;
if(cycle==2600)RxD<=1;
if(cycle==2700)RxD<=1;
if(cycle==2800)RxD<=1;
if(cycle==2900)RxD<=0;
if(cycle==3000)RxD<=1;
if(cycle==3100)RxD<=1;
if(cycle==3200)RxD<=0;
if(cycle==3300)RxD<=0;
if(cycle==3400)RxD<=1;
if(cycle==3500)RxD<=1;
if(cycle==3600)RxD<=1;
if(cycle==3700)RxD<=0;
if(cycle==3800)RxD<=0;
if(cycle==3900)RxD<=1;
if(cycle==4000)RxD<=0;
if(cycle==4100)RxD<=1;
if(cycle==4200)RxD<=0;
if(cycle==4300)RxD<=1;
if(cycle==4400)RxD<=0;
if(cycle==4500)RxD<=0;
if(cycle==4600)RxD<=1;
if(cycle==4700)RxD<=0;
if(cycle==4800)RxD<=0;
if(cycle==4900)RxD<=1;
if(cycle==5000)RxD<=1;
if(cycle==5100)RxD<=1;
if(cycle==5200)RxD<=0;
if(cycle==5300)RxD<=0;
if(cycle==5400)RxD<=0;
if(cycle==5500)RxD<=0;
if(cycle==5600)RxD<=1;
if(cycle==5700)RxD<=1;
if(cycle==5800)RxD<=0;
if(cycle==5900)RxD<=0;
if(cycle==6000)RxD<=1;
if(cycle==6100)RxD<=1;
if(cycle==6200)RxD<=0;
if(cycle==6300)RxD<=0;
if(cycle==6400)RxD<=1;
if(cycle==6500)RxD<=1;
if(cycle==6600)RxD<=0;
if(cycle==6700)RxD<=1;
if(cycle==6800)RxD<=1;
if(cycle==6900)RxD<=1;
if(cycle==7000)RxD<=0;
if(cycle==7100)RxD<=1;
if(cycle==7200)RxD<=0;
if(cycle==7300)RxD<=1;
if(cycle==7400)RxD<=1;
if(cycle==7500)RxD<=1;
if(cycle==7600)RxD<=1;
if(cycle==7700)RxD<=1;
if(cycle==7800)RxD<=1;
if(cycle==7900)RxD<=0;
if(cycle==8000)RxD<=1;
if(cycle==8100)RxD<=1;
if(cycle==8200)RxD<=0;
if(cycle==8300)RxD<=1;
if(cycle==8400)RxD<=1;
if(cycle==8500)RxD<=0;
if(cycle==8600)RxD<=1;
if(cycle==8700)RxD<=0;
if(cycle==8800)RxD<=0;
if(cycle==8900)RxD<=1;
if(cycle==9000)RxD<=0;
if(cycle==9100)RxD<=1;
if(cycle==9200)RxD<=0;
if(cycle==9300)RxD<=0;
if(cycle==9400)RxD<=1;
if(cycle==9500)RxD<=1;
if(cycle==9600)RxD<=1;
if(cycle==9700)RxD<=1;
if(cycle==9800)RxD<=1;
if(cycle==9900)RxD<=1;
if(cycle==10000)RxD<=1;
if(cycle==10100)RxD<=1;
if(cycle==10200)RxD<=0;
if(cycle==10300)RxD<=0;
if(cycle==10400)RxD<=0;
if(cycle==10500)RxD<=0;
if(cycle==10600)RxD<=1;
if(cycle==10700)RxD<=0;
if(cycle==10800)RxD<=0;
if(cycle==10900)RxD<=0;
if(cycle==11000)RxD<=0;
if(cycle==11100)RxD<=1;
if(cycle==11200)RxD<=0;
if(cycle==11300)RxD<=0;
if(cycle==11400)RxD<=0;
if(cycle==11500)RxD<=0;
if(cycle==11600)RxD<=0;
if(cycle==11700)RxD<=0;
if(cycle==11800)RxD<=1;
if(cycle==11900)RxD<=1;
if(cycle==12000)RxD<=0;
if(cycle==12100)RxD<=1;
if(cycle==12200)RxD<=0;
if(cycle==12300)RxD<=0;
if(cycle==12400)RxD<=1;
if(cycle==12500)RxD<=0;
if(cycle==12600)RxD<=0;
if(cycle==12700)RxD<=0;
if(cycle==12800)RxD<=0;
if(cycle==12900)RxD<=0;
if(cycle==13000)RxD<=1;
if(cycle==13100)RxD<=1;
if(cycle==13200)RxD<=0;
if(cycle==13300)RxD<=0;
if(cycle==13400)RxD<=0;
if(cycle==13500)RxD<=1;
if(cycle==13600)RxD<=0;
if(cycle==13700)RxD<=1;
if(cycle==13800)RxD<=1;
if(cycle==13900)RxD<=0;
if(cycle==14000)RxD<=1;
if(cycle==14100)RxD<=1;
if(cycle==14200)RxD<=0;
if(cycle==14300)RxD<=0;
if(cycle==14400)RxD<=0;
if(cycle==14500)RxD<=0;
if(cycle==14600)RxD<=0;
if(cycle==14700)RxD<=0;
if(cycle==14800)RxD<=0;
if(cycle==14900)RxD<=0;
if(cycle==15000)RxD<=0;
if(cycle==15100)RxD<=1;
if(cycle==15200)RxD<=0;
if(cycle==15300)RxD<=1;
if(cycle==15400)RxD<=0;
if(cycle==15500)RxD<=1;
if(cycle==15600)RxD<=0;
if(cycle==15700)RxD<=0;
if(cycle==15800)RxD<=1;
if(cycle==15900)RxD<=0;
if(cycle==16000)RxD<=0;
if(cycle==16100)RxD<=1;
if(cycle==16200)RxD<=0;
if(cycle==16300)RxD<=1;
if(cycle==16400)RxD<=0;
if(cycle==16500)RxD<=1;
if(cycle==16600)RxD<=1;
if(cycle==16700)RxD<=0;
if(cycle==16800)RxD<=0;
if(cycle==16900)RxD<=1;
if(cycle==17000)RxD<=0;
if(cycle==17100)RxD<=1;
if(cycle==17200)RxD<=0;
if(cycle==17300)RxD<=0;
if(cycle==17400)RxD<=1;
if(cycle==17500)RxD<=1;
if(cycle==17600)RxD<=0;
if(cycle==17700)RxD<=1;
if(cycle==17800)RxD<=1;
if(cycle==17900)RxD<=1;
if(cycle==18000)RxD<=1;
if(cycle==18100)RxD<=1;
if(cycle==18200)RxD<=0;
if(cycle==18300)RxD<=1;
if(cycle==18400)RxD<=1;
if(cycle==18500)RxD<=0;
if(cycle==18600)RxD<=0;
if(cycle==18700)RxD<=0;
if(cycle==18800)RxD<=0;
if(cycle==18900)RxD<=1;
if(cycle==19000)RxD<=1;
if(cycle==19100)RxD<=1;
if(cycle==19200)RxD<=0;
if(cycle==19300)RxD<=0;
if(cycle==19400)RxD<=1;
if(cycle==19500)RxD<=1;
if(cycle==19600)RxD<=0;
if(cycle==19700)RxD<=1;
if(cycle==19800)RxD<=0;
if(cycle==19900)RxD<=1;
if(cycle==20000)RxD<=0;
if(cycle==20100)RxD<=1;
if(cycle==20200)RxD<=0;
if(cycle==20300)RxD<=1;
if(cycle==20400)RxD<=0;
if(cycle==20500)RxD<=1;
if(cycle==20600)RxD<=0;
if(cycle==20700)RxD<=0;
if(cycle==20800)RxD<=0;
if(cycle==20900)RxD<=1;
if(cycle==21000)RxD<=0;
if(cycle==21100)RxD<=1;
if(cycle==21200)RxD<=0;
if(cycle==21300)RxD<=0;
if(cycle==21400)RxD<=0;
if(cycle==21500)RxD<=1;
if(cycle==21600)RxD<=0;
if(cycle==21700)RxD<=1;
if(cycle==21800)RxD<=0;
if(cycle==21900)RxD<=0;
if(cycle==22000)RxD<=0;
if(cycle==22100)RxD<=1;
if(cycle==22200)RxD<=0;
if(cycle==22300)RxD<=1;
if(cycle==22400)RxD<=0;
if(cycle==22500)RxD<=0;
if(cycle==22600)RxD<=0;
if(cycle==22700)RxD<=1;
if(cycle==22800)RxD<=1;
if(cycle==22900)RxD<=1;
if(cycle==23000)RxD<=0;
if(cycle==23100)RxD<=1;
if(cycle==23200)RxD<=0;
if(cycle==23300)RxD<=1;
if(cycle==23400)RxD<=1;
if(cycle==23500)RxD<=0;
if(cycle==23600)RxD<=0;
if(cycle==23700)RxD<=1;
if(cycle==23800)RxD<=0;
if(cycle==23900)RxD<=0;
if(cycle==24000)RxD<=0;
if(cycle==24100)RxD<=1;
if(cycle==24200)RxD<=0;
if(cycle==24300)RxD<=0;
if(cycle==24400)RxD<=1;
if(cycle==24500)RxD<=0;
if(cycle==24600)RxD<=1;
if(cycle==24700)RxD<=1;
if(cycle==24800)RxD<=0;
if(cycle==24900)RxD<=0;
if(cycle==25000)RxD<=1;
if(cycle==25100)RxD<=1;
if(cycle==25200)RxD<=0;
if(cycle==25300)RxD<=0;
if(cycle==25400)RxD<=1;
if(cycle==25500)RxD<=0;
if(cycle==25600)RxD<=1;
if(cycle==25700)RxD<=1;
if(cycle==25800)RxD<=1;
if(cycle==25900)RxD<=0;
if(cycle==26000)RxD<=0;
if(cycle==26100)RxD<=1;
if(cycle==26200)RxD<=0;
if(cycle==26300)RxD<=0;
if(cycle==26400)RxD<=1;
if(cycle==26500)RxD<=0;
if(cycle==26600)RxD<=1;
if(cycle==26700)RxD<=1;
if(cycle==26800)RxD<=1;
if(cycle==26900)RxD<=1;
if(cycle==27000)RxD<=1;
if(cycle==27100)RxD<=1;
if(cycle==27200)RxD<=0;
if(cycle==27300)RxD<=1;
if(cycle==27400)RxD<=0;
if(cycle==27500)RxD<=0;
if(cycle==27600)RxD<=0;
if(cycle==27700)RxD<=1;
if(cycle==27800)RxD<=1;
if(cycle==27900)RxD<=1;
if(cycle==28000)RxD<=0;
if(cycle==28100)RxD<=1;
if(cycle==28200)RxD<=0;
if(cycle==28300)RxD<=0;
if(cycle==28400)RxD<=0;
if(cycle==28500)RxD<=1;
if(cycle==28600)RxD<=0;
if(cycle==28700)RxD<=0;
if(cycle==28800)RxD<=1;
if(cycle==28900)RxD<=1;
if(cycle==29000)RxD<=1;
if(cycle==29100)RxD<=1;
if(cycle==29200)RxD<=0;
if(cycle==29300)RxD<=1;
if(cycle==29400)RxD<=1;
if(cycle==29500)RxD<=1;
if(cycle==29600)RxD<=1;
if(cycle==29700)RxD<=0;
if(cycle==29800)RxD<=0;
if(cycle==29900)RxD<=0;
if(cycle==30000)RxD<=1;
if(cycle==30100)RxD<=1;
if(cycle==30200)RxD<=0;
if(cycle==30300)RxD<=0;
if(cycle==30400)RxD<=0;
if(cycle==30500)RxD<=1;
if(cycle==30600)RxD<=0;
if(cycle==30700)RxD<=1;
if(cycle==30800)RxD<=0;
if(cycle==30900)RxD<=1;
if(cycle==31000)RxD<=0;
if(cycle==31100)RxD<=1;
if(cycle==31200)RxD<=0;
if(cycle==31300)RxD<=0;
if(cycle==31400)RxD<=1;
if(cycle==31500)RxD<=0;
if(cycle==31600)RxD<=1;
if(cycle==31700)RxD<=0;
if(cycle==31800)RxD<=0;
if(cycle==31900)RxD<=1;
if(cycle==32000)RxD<=0;
if(cycle==32100)RxD<=1;
if(cycle==32200)RxD<=0;
if(cycle==32300)RxD<=0;
if(cycle==32400)RxD<=0;
if(cycle==32500)RxD<=0;
if(cycle==32600)RxD<=0;
if(cycle==32700)RxD<=0;
if(cycle==32800)RxD<=0;
if(cycle==32900)RxD<=0;
if(cycle==33000)RxD<=0;
if(cycle==33100)RxD<=1;
if(cycle==33200)RxD<=0;
if(cycle==33300)RxD<=0;
if(cycle==33400)RxD<=0;
if(cycle==33500)RxD<=0;
if(cycle==33600)RxD<=0;
if(cycle==33700)RxD<=0;
if(cycle==33800)RxD<=0;
if(cycle==33900)RxD<=0;
if(cycle==34000)RxD<=0;
if(cycle==34100)RxD<=1;
if(cycle==34200)RxD<=0;
if(cycle==34300)RxD<=0;
if(cycle==34400)RxD<=0;
if(cycle==34500)RxD<=0;
if(cycle==34600)RxD<=0;
if(cycle==34700)RxD<=0;
if(cycle==34800)RxD<=0;
if(cycle==34900)RxD<=0;
if(cycle==35000)RxD<=0;
if(cycle==35100)RxD<=1;
if(cycle==35200)RxD<=0;
if(cycle==35300)RxD<=0;
if(cycle==35400)RxD<=0;
if(cycle==35500)RxD<=0;
if(cycle==35600)RxD<=0;
if(cycle==35700)RxD<=0;
if(cycle==35800)RxD<=0;
if(cycle==35900)RxD<=0;
if(cycle==36000)RxD<=0;
if(cycle==36100)RxD<=1;
if(cycle==36200)RxD<=0;
if(cycle==36300)RxD<=0;
if(cycle==36400)RxD<=0;
if(cycle==36500)RxD<=0;
if(cycle==36600)RxD<=0;
if(cycle==36700)RxD<=0;
if(cycle==36800)RxD<=0;
if(cycle==36900)RxD<=0;
if(cycle==37000)RxD<=0;
if(cycle==37100)RxD<=1;
if(cycle==37200)RxD<=0;
if(cycle==37300)RxD<=0;
if(cycle==37400)RxD<=0;
if(cycle==37500)RxD<=0;
if(cycle==37600)RxD<=0;
if(cycle==37700)RxD<=0;
if(cycle==37800)RxD<=0;
if(cycle==37900)RxD<=0;
if(cycle==38000)RxD<=0;
if(cycle==38100)RxD<=1;
if(cycle==38200)RxD<=0;
if(cycle==38300)RxD<=0;
if(cycle==38400)RxD<=0;
if(cycle==38500)RxD<=0;
if(cycle==38600)RxD<=0;
if(cycle==38700)RxD<=0;
if(cycle==38800)RxD<=0;
if(cycle==38900)RxD<=0;
if(cycle==39000)RxD<=0;
if(cycle==39100)RxD<=1;
if(cycle==39200)RxD<=0;
if(cycle==39300)RxD<=0;
if(cycle==39400)RxD<=0;
if(cycle==39500)RxD<=0;
if(cycle==39600)RxD<=0;
if(cycle==39700)RxD<=0;
if(cycle==39800)RxD<=0;
if(cycle==39900)RxD<=0;
if(cycle==40000)RxD<=0;
if(cycle==40100)RxD<=1;
if(cycle==40200)RxD<=0;
if(cycle==40300)RxD<=0;
if(cycle==40400)RxD<=0;
if(cycle==40500)RxD<=0;
if(cycle==40600)RxD<=0;
if(cycle==40700)RxD<=0;
if(cycle==40800)RxD<=0;
if(cycle==40900)RxD<=0;
if(cycle==41000)RxD<=0;
if(cycle==41100)RxD<=1;
if(cycle==41200)RxD<=0;
if(cycle==41300)RxD<=0;
if(cycle==41400)RxD<=0;
if(cycle==41500)RxD<=0;
if(cycle==41600)RxD<=0;
if(cycle==41700)RxD<=0;
if(cycle==41800)RxD<=0;
if(cycle==41900)RxD<=0;
if(cycle==42000)RxD<=0;
if(cycle==42100)RxD<=1;
if(cycle==42200)RxD<=0;
if(cycle==42300)RxD<=0;
if(cycle==42400)RxD<=0;
if(cycle==42500)RxD<=0;
if(cycle==42600)RxD<=0;
if(cycle==42700)RxD<=0;
if(cycle==42800)RxD<=0;
if(cycle==42900)RxD<=0;
if(cycle==43000)RxD<=0;
if(cycle==43100)RxD<=1;
if(cycle==43200)RxD<=0;
if(cycle==43300)RxD<=0;
if(cycle==43400)RxD<=0;
if(cycle==43500)RxD<=0;
if(cycle==43600)RxD<=0;
if(cycle==43700)RxD<=0;
if(cycle==43800)RxD<=0;
if(cycle==43900)RxD<=0;
if(cycle==44000)RxD<=0;
if(cycle==44100)RxD<=1;
if(cycle==44200)RxD<=0;
if(cycle==44300)RxD<=0;
if(cycle==44400)RxD<=0;
if(cycle==44500)RxD<=0;
if(cycle==44600)RxD<=0;
if(cycle==44700)RxD<=0;
if(cycle==44800)RxD<=0;
if(cycle==44900)RxD<=0;
if(cycle==45000)RxD<=0;
if(cycle==45100)RxD<=1;
if(cycle==45200)RxD<=0;
if(cycle==45300)RxD<=0;
if(cycle==45400)RxD<=0;
if(cycle==45500)RxD<=0;
if(cycle==45600)RxD<=0;
if(cycle==45700)RxD<=0;
if(cycle==45800)RxD<=0;
if(cycle==45900)RxD<=0;
if(cycle==46000)RxD<=0;
if(cycle==46100)RxD<=1;
if(cycle==46200)RxD<=0;
if(cycle==46300)RxD<=0;
if(cycle==46400)RxD<=0;
if(cycle==46500)RxD<=0;
if(cycle==46600)RxD<=0;
if(cycle==46700)RxD<=0;
if(cycle==46800)RxD<=0;
if(cycle==46900)RxD<=0;
if(cycle==47000)RxD<=0;
if(cycle==47100)RxD<=1;
if(cycle==47200)RxD<=0;
if(cycle==47300)RxD<=0;
if(cycle==47400)RxD<=0;
if(cycle==47500)RxD<=0;
if(cycle==47600)RxD<=0;
if(cycle==47700)RxD<=0;
if(cycle==47800)RxD<=0;
if(cycle==47900)RxD<=0;
if(cycle==48000)RxD<=0;
if(cycle==48100)RxD<=1;
if(cycle==48200)RxD<=0;
if(cycle==48300)RxD<=0;
if(cycle==48400)RxD<=0;
if(cycle==48500)RxD<=0;
if(cycle==48600)RxD<=0;
if(cycle==48700)RxD<=0;
if(cycle==48800)RxD<=0;
if(cycle==48900)RxD<=0;
if(cycle==49000)RxD<=0;
if(cycle==49100)RxD<=1;
if(cycle==49200)RxD<=0;
if(cycle==49300)RxD<=0;
if(cycle==49400)RxD<=0;
if(cycle==49500)RxD<=0;
if(cycle==49600)RxD<=0;
if(cycle==49700)RxD<=0;
if(cycle==49800)RxD<=0;
if(cycle==49900)RxD<=0;
if(cycle==50000)RxD<=0;
if(cycle==50100)RxD<=1;
if(cycle==50200)RxD<=0;
if(cycle==50300)RxD<=0;
if(cycle==50400)RxD<=0;
if(cycle==50500)RxD<=0;
if(cycle==50600)RxD<=0;
if(cycle==50700)RxD<=0;
if(cycle==50800)RxD<=0;
if(cycle==50900)RxD<=0;
if(cycle==51000)RxD<=0;
if(cycle==51100)RxD<=1;
if(cycle==51200)RxD<=0;
if(cycle==51300)RxD<=0;
if(cycle==51400)RxD<=0;
if(cycle==51500)RxD<=0;
if(cycle==51600)RxD<=0;
if(cycle==51700)RxD<=0;
if(cycle==51800)RxD<=0;
if(cycle==51900)RxD<=0;
if(cycle==52000)RxD<=0;
if(cycle==52100)RxD<=1;
if(cycle==52200)RxD<=0;
if(cycle==52300)RxD<=1;
if(cycle==52400)RxD<=1;
if(cycle==52500)RxD<=1;
if(cycle==52600)RxD<=0;
if(cycle==52700)RxD<=0;
if(cycle==52800)RxD<=0;
if(cycle==52900)RxD<=0;
if(cycle==53000)RxD<=1;
if(cycle==53100)RxD<=1;
if(cycle==53200)RxD<=0;
if(cycle==53300)RxD<=0;
if(cycle==53400)RxD<=1;
if(cycle==53500)RxD<=0;
if(cycle==53600)RxD<=0;
if(cycle==53700)RxD<=1;
if(cycle==53800)RxD<=1;
if(cycle==53900)RxD<=0;
if(cycle==54000)RxD<=0;
if(cycle==54100)RxD<=1;
if(cycle==54200)RxD<=0;
if(cycle==54300)RxD<=1;
if(cycle==54400)RxD<=1;
if(cycle==54500)RxD<=0;
if(cycle==54600)RxD<=1;
if(cycle==54700)RxD<=0;
if(cycle==54800)RxD<=0;
if(cycle==54900)RxD<=0;
if(cycle==55000)RxD<=0;
if(cycle==55100)RxD<=1;
if(cycle==55200)RxD<=0;
if(cycle==55300)RxD<=0;
if(cycle==55400)RxD<=1;
if(cycle==55500)RxD<=0;
if(cycle==55600)RxD<=1;
if(cycle==55700)RxD<=1;
if(cycle==55800)RxD<=0;
if(cycle==55900)RxD<=0;
if(cycle==56000)RxD<=0;
if(cycle==56100)RxD<=1;
if(cycle==56200)RxD<=0;
if(cycle==56300)RxD<=0;
if(cycle==56400)RxD<=0;
if(cycle==56500)RxD<=1;
if(cycle==56600)RxD<=0;
if(cycle==56700)RxD<=1;
if(cycle==56800)RxD<=0;
if(cycle==56900)RxD<=0;
if(cycle==57000)RxD<=0;
if(cycle==57100)RxD<=1;
if(cycle==57200)RxD<=0;
if(cycle==57300)RxD<=0;
if(cycle==57400)RxD<=1;
if(cycle==57500)RxD<=1;
if(cycle==57600)RxD<=0;
if(cycle==57700)RxD<=0;
if(cycle==57800)RxD<=1;
if(cycle==57900)RxD<=0;
if(cycle==58000)RxD<=0;
if(cycle==58100)RxD<=1;
if(cycle==58200)RxD<=0;
if(cycle==58300)RxD<=1;
if(cycle==58400)RxD<=1;
if(cycle==58500)RxD<=1;
if(cycle==58600)RxD<=0;
if(cycle==58700)RxD<=0;
if(cycle==58800)RxD<=1;
if(cycle==58900)RxD<=1;
if(cycle==59000)RxD<=0;
if(cycle==59100)RxD<=1;
if(cycle==59200)RxD<=0;
if(cycle==59300)RxD<=1;
if(cycle==59400)RxD<=1;
if(cycle==59500)RxD<=1;
if(cycle==59600)RxD<=1;
if(cycle==59700)RxD<=0;
if(cycle==59800)RxD<=0;
if(cycle==59900)RxD<=1;
if(cycle==60000)RxD<=0;
if(cycle==60100)RxD<=1;
if(cycle==60200)RxD<=0;
if(cycle==60300)RxD<=1;
if(cycle==60400)RxD<=1;
if(cycle==60500)RxD<=1;
if(cycle==60600)RxD<=1;
if(cycle==60700)RxD<=0;
if(cycle==60800)RxD<=1;
if(cycle==60900)RxD<=0;
if(cycle==61000)RxD<=0;
if(cycle==61100)RxD<=1;
if(cycle==61200)RxD<=0;
if(cycle==61300)RxD<=1;
if(cycle==61400)RxD<=1;
if(cycle==61500)RxD<=1;
if(cycle==61600)RxD<=0;
if(cycle==61700)RxD<=0;
if(cycle==61800)RxD<=1;
if(cycle==61900)RxD<=0;
if(cycle==62000)RxD<=1;
if(cycle==62100)RxD<=1;
if(cycle==62200)RxD<=0;
if(cycle==62300)RxD<=0;
if(cycle==62400)RxD<=1;
if(cycle==62500)RxD<=0;
if(cycle==62600)RxD<=0;
if(cycle==62700)RxD<=0;
if(cycle==62800)RxD<=1;
if(cycle==62900)RxD<=0;
if(cycle==63000)RxD<=0;
if(cycle==63100)RxD<=1;
if(cycle==63200)RxD<=0;
if(cycle==63300)RxD<=0;
if(cycle==63400)RxD<=1;
if(cycle==63500)RxD<=1;
if(cycle==63600)RxD<=1;
if(cycle==63700)RxD<=0;
if(cycle==63800)RxD<=0;
if(cycle==63900)RxD<=1;
if(cycle==64000)RxD<=1;
if(cycle==64100)RxD<=1;
			
			
		end
	end


	always @ (posedge clk)
	begin
		cycle <= cycle + 32'd1;
	end

endmodule

